module test_bench();
	
	reg valid;
	reg [31:0]x0;
	reg [31:0]y0;
	reg [31:0]z0;
	reg [31:0]n;
	wire [31:0]x;
	wire [31:0]y;
	wire [31:0]z;

	initial
		begin
			
		end


endmodule